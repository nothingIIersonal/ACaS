library verilog;
use verilog.vl_types.all;
entity lab42_vlg_vec_tst is
end lab42_vlg_vec_tst;
