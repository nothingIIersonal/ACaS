library verilog;
use verilog.vl_types.all;
entity lab12_vlg_vec_tst is
end lab12_vlg_vec_tst;
