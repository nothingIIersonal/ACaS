library verilog;
use verilog.vl_types.all;
entity lab21_vlg_vec_tst is
end lab21_vlg_vec_tst;
