library verilog;
use verilog.vl_types.all;
entity lab22_vlg_vec_tst is
end lab22_vlg_vec_tst;
