library verilog;
use verilog.vl_types.all;
entity lab23_vlg_vec_tst is
end lab23_vlg_vec_tst;
