library verilog;
use verilog.vl_types.all;
entity lab41_vlg_vec_tst is
end lab41_vlg_vec_tst;
