library verilog;
use verilog.vl_types.all;
entity lab21_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab21_vlg_check_tst;
