library verilog;
use verilog.vl_types.all;
entity lab21 is
    port(
        F               : out    vl_logic;
        D0              : in     vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        D2              : in     vl_logic;
        D1              : in     vl_logic;
        D3              : in     vl_logic;
        D5              : in     vl_logic;
        D4              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic
    );
end lab21;
